module pwm_test(CLOCK_50,SW,KEY,LEDG);
paramter WIDTH = 12;
input wire CLOCK_50;
input wire[17:0] SW;
input wire[3:0] KEY;
output wire[8:0] LEDG;
wire[WIDTH-1:0] 
endmodule
